LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY dadda_16x16_multiplier is
PORT(A,B: IN std_logic_vector(15 downto 0);
     M: OUT std_logic_vector(31 downto 0));

END dadda_16x16_multiplier;


ARCHITECTURE a1 of dadda_16x16_multiplier is


COMPONENT FULLADD is
PORT(A,B,C: IN std_logic;
     Sum,Cout: OUT std_logic);

END COMPONENT;

COMPONENT HALFADD is
PORT(A,B: IN std_logic;
     Sum,Cout: OUT std_logic);

END COMPONENT;

COMPONENT brentkung_32bit_adder is
PORT ( A,B : IN STD_LOGIC_VECTOR(31 downto 0) ;
       Cin: IN std_logic; 
       Sum : OUT STD_LOGIC_VECTOR(31 downto 0)  ;
       Cout: OUT std_logic);

END COMPONENT; 

--    signals

signal nocarry: std_logic;
signal Ain,Bin: std_logic_vector(31 downto 0);

-- some dummy signals

signal dum0,dum1,dum2,dum3,dum4,dum5,dum6,dum7,dum8,dum9,dum10,dum11,dum12,dum13,dum14,dum15,dum16,dum17,dum18,dum19,dum20,dum21,dum22,dum23,dum24,dum25,dum26,dum27,dum28,dum29,dum30: STD_LOGIC;

signal dum31,dum32,dum33,dum34,dum35,dum36,dum37,dum38,dum39,dum40,dum41,dum42,dum43,dum44,dum45,dum46,dum47,dum48,dum49,dum50,dum51,dum52,dum53,dum54,dum55,dum56,dum57,dum58,dum59,dum60: STD_LOGIC;

signal dum61,dum62,dum63,dum64,dum65,dum66,dum67,dum68,dum69,dum70,dum71,dum72,dum73,dum74,dum75,dum76,dum77,dum78,dum79,dum80,dum81,dum82,dum83,dum84,dum85,dum86,dum87,dum88,dum89,dum90: STD_LOGIC;

signal dum91,dum92,dum93,dum94,dum95,dum96,dum97,dum98,dum99,dum100: STD_LOGIC;

signal dum101,dum102,dum103,dum104,dum105,dum106,dum107,dum108,dum109,dum110,dum111,dum112,dum113,dum114,dum115,dum116,dum117,dum118,dum119,dum120,dum121,dum122,dum123,dum124,dum125,dum126,dum127,dum128,dum129,dum130: STD_LOGIC;

signal dum131,dum132,dum133,dum134,dum135,dum136,dum137,dum138,dum139,dum140,dum141,dum142,dum143,dum144,dum145,dum146,dum147,dum148,dum149,dum150,dum151,dum152,dum153,dum154,dum155,dum156,dum157,dum158,dum159,dum160: STD_LOGIC;

signal dum161,dum162,dum163,dum164,dum165,dum166,dum167,dum168,dum169,dum170,dum171,dum172,dum173,dum174,dum175,dum176,dum177,dum178,dum179,dum180,dum181,dum182,dum183,dum184,dum185,dum186,dum187,dum188,dum189,dum190: STD_LOGIC;

signal dum191,dum192,dum193,dum194,dum195,dum196,dum197,dum198,dum199,dum200: STD_LOGIC;

signal dum201,dum202,dum203,dum204,dum205,dum206,dum207,dum208,dum209,dum210,dum211,dum212,dum213,dum214,dum215,dum216,dum217,dum218,dum219,dum220,dum221,dum222,dum223,dum224,dum225,dum226,dum227,dum228,dum229,dum230: STD_LOGIC;

signal dum231,dum232,dum233,dum234,dum235,dum236,dum237,dum238,dum239,dum240,dum241,dum242,dum243,dum244,dum245,dum246,dum247,dum248,dum249,dum250,dum251,dum252,dum253,dum254,dum255: STD_LOGIC;

--starting signals name

signal A0B0,A0B1,A1B0,A0B2,A1B1,A2B0,A0B3,A1B2,A2B1,A3B0,A0B4,A1B3,A2B2,A3B1,A4B0,A0B5,A1B4,A2B3,A3B2,A4B1,A5B0,A0B6,A1B5,A2B4,A3B3,A4B2,A5B1,A6B0,A0B7,A1B6,A2B5,A3B4,A4B3,A5B2,A6B1,A7B0,A0B8,A1B7,A2B6,A3B5,A4B4,A5B3,A6B2,A7B1,A8B0,A0B9,A1B8,A2B7,A3B6,A4B5,A5B4,A6B3,A7B2,A8B1,A9B0,A0B10,A1B9,A2B8,A3B7,A4B6,A5B5,A6B4,A7B3,A8B2,A9B1,A10B0,A0B11,A1B10,A2B9,A3B8,A4B7,A5B6,A6B5,A7B4,A8B3,A9B2,A10B1,A11B0,A0B12,A1B11,A2B10,A3B9,A4B8,A5B7,A6B6,A7B5,A8B4,A9B3,A10B2,A11B1,A12B0,A0B13,A1B12,A2B11,A3B10,A4B9,A5B8,A6B7,A7B6,A8B5,A9B4,A10B3,A11B2,A12B1,A13B0: std_logic;
signal A0B14,A1B13,A2B12,A3B11,A4B10,A5B9,A6B8,A7B7,A8B6,A9B5,A10B4,A11B3,A12B2,A13B1,A14B0,A0B15,A1B14,A2B13,A3B12,A4B11,A5B10,A6B9,A7B8,A8B7,A9B6,A10B5,A11B4,A12B3,A13B2,A14B1,A15B0,A1B15,A2B14,A3B13,A4B12,A5B11,A6B10,A7B9,A8B8,A9B7,A10B6,A11B5,A12B4,A13B3,A14B2,A15B1,A2B15,A3B14,A4B13,A5B12,A6B11,A7B10,A8B9,A9B8,A10B7,A11B6,A12B5,A13B4,A14B3,A15B2,A3B15,A4B14,A5B13,A6B12,A7B11,A8B10,A9B9,A10B8,A11B7,A12B6,A13B5,A14B4,A15B3,A4B15,A5B14,A6B13,A7B12,A8B11,A9B10,A10B9,A11B8,A12B7,A13B6,A14B5,A15B4: std_logic;
signal A5B15,A6B14,A7B13,A8B12,A9B11,A10B10,A11B9,A12B8,A13B7,A14B6,A15B5,A6B15,A7B14,A8B13,A9B12,A10B11,A11B10,A12B9,A13B8,A14B7,A15B6,A7B15,A8B14,A9B13,A10B12,A11B11,A12B10,A13B9,A14B8,A15B7,A8B15,A9B14,A10B13,A11B12,A12B11,A13B10,A14B9,A15B8,A9B15,A10B14,A11B13,A12B12,A13B11,A14B10,A15B9: std_logic;
signal A10B15,A11B14,A12B13,A13B12,A14B11,A15B10,A11B15,A12B14,A13B13,A14B12,A15B11,A12B15,A13B14,A14B13,A15B12,A13B15,A14B14,A15B13,A14B15,A15B14,A15B15: std_logic;


--some signals which will be used in further operation

signal Sn1L1_14_Sn2L1_1,Sn1L1_15_Sn2L1_1,Sn1L1_16_Sn2L1_1,Sn1L1_17_Sn2L1_1,Sn1L1_18_Sn2L1_1,Sn1L1_19_Sn2L1_1:std_logic;
signal Sn1L1_15_Sn2L1_2,Sn1L1_16_Sn2L1_2,Sn1L1_17_Sn2L1_2,Sn1L1_18_Sn2L1_2,Sn1L1_19_Sn2L1_2,Sn1L1_20_Sn2L1_2:std_logic;
signal Sn1L1_15_Sn2L1_3,Sn1L1_16_Sn2L1_3,Sn1L1_17_Sn2L1_3,Sn1L1_18_Sn2L1_3:std_logic;
signal Sn1L1_16_Sn2L1_4,Sn1L1_17_Sn2L1_4,Sn1L1_18_Sn2L1_4,Sn1L1_19_Sn2L1_4:std_logic;
signal Sn1L1_16_Sn2L1_5,Sn1L1_17_Sn2L1_5:std_logic;
signal Sn1L1_17_Sn2L1_6,Sn1L1_18_Sn2L1_6:std_logic;
signal Sn1L2_10_Sn2L2_1,Sn1L2_11_Sn2L2_1,Sn1L2_12_Sn2L2_1,Sn1L2_13_Sn2L2_1,Sn1L2_14_Sn2L2_1,Sn1L2_15_Sn2L2_1,Sn1L2_16_Sn2L2_1,Sn1L2_17_Sn2L2_1,Sn1L2_18_Sn2L2_1,Sn1L2_19_Sn2L2_1,Sn1L2_20_Sn2L2_1,Sn1L2_21_Sn2L2_1,Sn1L2_22_Sn2L2_1,Sn1L2_23_Sn2L2_1:std_logic;
signal Sn1L2_11_Sn2L2_2,Sn1L2_12_Sn2L2_2,Sn1L2_13_Sn2L2_2,Sn1L2_14_Sn2L2_2,Sn1L2_15_Sn2L2_2,Sn1L2_16_Sn2L2_2,Sn1L2_17_Sn2L2_2,Sn1L2_18_Sn2L2_2,Sn1L2_19_Sn2L2_2,Sn1L2_20_Sn2L2_2,Sn1L2_21_Sn2L2_2,Sn1L2_22_Sn2L2_2,Sn1L2_23_Sn2L2_2,Sn1L2_24_Sn2L2_2:std_logic;
signal Sn1L2_11_Sn2L2_3,Sn1L2_12_Sn2L2_3,Sn1L2_13_Sn2L2_3,Sn1L2_14_Sn2L2_3,Sn1L2_15_Sn2L2_3,Sn1L2_16_Sn2L2_3,Sn1L2_17_Sn2L2_3,Sn1L2_18_Sn2L2_3,Sn1L2_19_Sn2L2_3,Sn1L2_20_Sn2L2_3,Sn1L2_21_Sn2L2_3,Sn1L2_22_Sn2L2_3:std_logic;
signal Sn1L2_12_Sn2L2_4,Sn1L2_13_Sn2L2_4,Sn1L2_14_Sn2L2_4,Sn1L2_15_Sn2L2_4,Sn1L2_16_Sn2L2_4,Sn1L2_17_Sn2L2_4,Sn1L2_18_Sn2L2_4,Sn1L2_19_Sn2L2_4,Sn1L2_20_Sn2L2_4,Sn1L2_21_Sn2L2_4,Sn1L2_22_Sn2L2_4,Sn1L2_23_Sn2L2_4:std_logic;
signal Sn1L2_12_Sn2L2_5,Sn1L2_13_Sn2L2_5,Sn1L2_14_Sn2L2_5,Sn1L2_15_Sn2L2_5,Sn1L2_16_Sn2L2_5,Sn1L2_17_Sn2L2_5,Sn1L2_18_Sn2L2_5,Sn1L2_19_Sn2L2_5,Sn1L2_20_Sn2L2_5,Sn1L2_21_Sn2L2_5:std_logic;
signal Sn1L2_13_Sn2L2_6,Sn1L2_14_Sn2L2_6,Sn1L2_15_Sn2L2_6,Sn1L2_16_Sn2L2_6,Sn1L2_17_Sn2L2_6,Sn1L2_18_Sn2L2_6,Sn1L2_19_Sn2L2_6,Sn1L2_20_Sn2L2_6,Sn1L2_21_Sn2L2_6,Sn1L2_22_Sn2L2_6:std_logic;
signal Sn1L2_13_Sn2L2_7,Sn1L2_14_Sn2L2_7,Sn1L2_15_Sn2L2_7,Sn1L2_16_Sn2L2_7,Sn1L2_17_Sn2L2_7,Sn1L2_18_Sn2L2_7,Sn1L2_19_Sn2L2_7,Sn1L2_20_Sn2L2_7:std_logic;
signal Sn1L2_14_Sn2L2_8,Sn1L2_15_Sn2L2_8,Sn1L2_16_Sn2L2_8,Sn1L2_17_Sn2L2_8,Sn1L2_18_Sn2L2_8,Sn1L2_19_Sn2L2_8,Sn1L2_20_Sn2L2_8,Sn1L2_21_Sn2L2_8:std_logic;
signal Sn1L3_7_Sn2L3_1,Sn1L3_8_Sn2L3_1,Sn1L3_9_Sn2L3_1,Sn1L3_10_Sn2L3_1,Sn1L3_11_Sn2L3_1,Sn1L3_12_Sn2L3_1,Sn1L3_13_Sn2L3_1,Sn1L3_14_Sn2L3_1,Sn1L3_15_Sn2L3_1,Sn1L3_16_Sn2L3_1,Sn1L3_17_Sn2L3_1,Sn1L3_18_Sn2L3_1,Sn1L3_19_Sn2L3_1,Sn1L3_20_Sn2L3_1,Sn1L3_21_Sn2L3_1,Sn1L3_22_Sn2L3_1,Sn1L3_23_Sn2L3_1,Sn1L3_24_Sn2L3_1,Sn1L3_25_Sn2L3_1,Sn1L3_26_Sn2L3_1:std_logic;
signal Sn1L3_8_Sn2L3_2,Sn1L3_9_Sn2L3_2,Sn1L3_10_Sn2L3_2,Sn1L3_11_Sn2L3_2,Sn1L3_12_Sn2L3_2,Sn1L3_13_Sn2L3_2,Sn1L3_14_Sn2L3_2,Sn1L3_15_Sn2L3_2,Sn1L3_16_Sn2L3_2,Sn1L3_17_Sn2L3_2,Sn1L3_18_Sn2L3_2,Sn1L3_19_Sn2L3_2,Sn1L3_20_Sn2L3_2,Sn1L3_21_Sn2L3_2,Sn1L3_22_Sn2L3_2,Sn1L3_23_Sn2L3_2,Sn1L3_24_Sn2L3_2,Sn1L3_25_Sn2L3_2,Sn1L3_26_Sn2L3_2,Sn1L3_27_Sn2L3_2:std_logic;
signal Sn1L3_8_Sn2L3_3,Sn1L3_9_Sn2L3_3,Sn1L3_10_Sn2L3_3,Sn1L3_11_Sn2L3_3,Sn1L3_12_Sn2L3_3,Sn1L3_13_Sn2L3_3,Sn1L3_14_Sn2L3_3,Sn1L3_15_Sn2L3_3,Sn1L3_16_Sn2L3_3,Sn1L3_17_Sn2L3_3,Sn1L3_18_Sn2L3_3,Sn1L3_19_Sn2L3_3,Sn1L3_20_Sn2L3_3,Sn1L3_21_Sn2L3_3,Sn1L3_22_Sn2L3_3,Sn1L3_23_Sn2L3_3,Sn1L3_24_Sn2L3_3,Sn1L3_25_Sn2L3_3:std_logic;
signal Sn1L3_9_Sn2L3_4,Sn1L3_10_Sn2L3_4,Sn1L3_11_Sn2L3_4,Sn1L3_12_Sn2L3_4,Sn1L3_13_Sn2L3_4,Sn1L3_14_Sn2L3_4,Sn1L3_15_Sn2L3_4,Sn1L3_16_Sn2L3_4,Sn1L3_17_Sn2L3_4,Sn1L3_18_Sn2L3_4,Sn1L3_19_Sn2L3_4,Sn1L3_20_Sn2L3_4,Sn1L3_21_Sn2L3_4,Sn1L3_22_Sn2L3_4,Sn1L3_23_Sn2L3_4,Sn1L3_24_Sn2L3_4,Sn1L3_25_Sn2L3_4,Sn1L3_26_Sn2L3_4:std_logic;
signal Sn1L3_9_Sn2L3_5,Sn1L3_10_Sn2L3_5,Sn1L3_11_Sn2L3_5,Sn1L3_12_Sn2L3_5,Sn1L3_13_Sn2L3_5,Sn1L3_14_Sn2L3_5,Sn1L3_15_Sn2L3_5,Sn1L3_16_Sn2L3_5,Sn1L3_17_Sn2L3_5,Sn1L3_18_Sn2L3_5,Sn1L3_19_Sn2L3_5,Sn1L3_20_Sn2L3_5,Sn1L3_21_Sn2L3_5,Sn1L3_22_Sn2L3_5,Sn1L3_23_Sn2L3_5,Sn1L3_24_Sn2L3_5:std_logic;
signal Sn1L3_10_Sn2L3_6,Sn1L3_11_Sn2L3_6,Sn1L3_12_Sn2L3_6,Sn1L3_13_Sn2L3_6,Sn1L3_14_Sn2L3_6,Sn1L3_15_Sn2L3_6,Sn1L3_16_Sn2L3_6,Sn1L3_17_Sn2L3_6,Sn1L3_18_Sn2L3_6,Sn1L3_19_Sn2L3_6,Sn1L3_20_Sn2L3_6,Sn1L3_21_Sn2L3_6,Sn1L3_22_Sn2L3_6,Sn1L3_23_Sn2L3_6,Sn1L3_24_Sn2L3_6,Sn1L3_25_Sn2L3_6:std_logic;
signal Sn1L4_5_Sn2L4_1,Sn1L4_6_Sn2L4_1,Sn1L4_7_Sn2L4_1,Sn1L4_8_Sn2L4_1,Sn1L4_9_Sn2L4_1,Sn1L4_10_Sn2L4_1,Sn1L4_11_Sn2L4_1,Sn1L4_12_Sn2L4_1,Sn1L4_13_Sn2L4_1,Sn1L4_14_Sn2L4_1,Sn1L4_15_Sn2L4_1,Sn1L4_16_Sn2L4_1,Sn1L4_17_Sn2L4_1,Sn1L4_18_Sn2L4_1,Sn1L4_19_Sn2L4_1,Sn1L4_20_Sn2L4_1,Sn1L4_21_Sn2L4_1,Sn1L4_22_Sn2L4_1,Sn1L4_23_Sn2L4_1,Sn1L4_24_Sn2L4_1,Sn1L4_25_Sn2L4_1,Sn1L4_26_Sn2L4_1,Sn1L4_27_Sn2L4_1,Sn1L4_28_Sn2L4_1: std_logic;
signal Sn1L4_6_Sn2L4_2,Sn1L4_7_Sn2L4_2,Sn1L4_8_Sn2L4_2,Sn1L4_9_Sn2L4_2,Sn1L4_10_Sn2L4_2,Sn1L4_11_Sn2L4_2,Sn1L4_12_Sn2L4_2,Sn1L4_13_Sn2L4_2,Sn1L4_14_Sn2L4_2,Sn1L4_15_Sn2L4_2,Sn1L4_16_Sn2L4_2,Sn1L4_17_Sn2L4_2,Sn1L4_18_Sn2L4_2,Sn1L4_19_Sn2L4_2,Sn1L4_20_Sn2L4_2,Sn1L4_21_Sn2L4_2,Sn1L4_22_Sn2L4_2,Sn1L4_23_Sn2L4_2,Sn1L4_24_Sn2L4_2,Sn1L4_25_Sn2L4_2,Sn1L4_26_Sn2L4_2,Sn1L4_27_Sn2L4_2,Sn1L4_28_Sn2L4_2,Sn1L4_29_Sn2L4_2: std_logic;
signal Sn1L4_6_Sn2L4_3,Sn1L4_7_Sn2L4_3,Sn1L4_8_Sn2L4_3,Sn1L4_9_Sn2L4_3,Sn1L4_10_Sn2L4_3,Sn1L4_11_Sn2L4_3,Sn1L4_12_Sn2L4_3,Sn1L4_13_Sn2L4_3,Sn1L4_14_Sn2L4_3,Sn1L4_15_Sn2L4_3,Sn1L4_16_Sn2L4_3,Sn1L4_17_Sn2L4_3,Sn1L4_18_Sn2L4_3,Sn1L4_19_Sn2L4_3,Sn1L4_20_Sn2L4_3,Sn1L4_21_Sn2L4_3,Sn1L4_22_Sn2L4_3,Sn1L4_23_Sn2L4_3,Sn1L4_24_Sn2L4_3,Sn1L4_25_Sn2L4_3,Sn1L4_26_Sn2L4_3,Sn1L4_27_Sn2L4_3: std_logic;
signal Sn1L4_7_Sn2L4_4,Sn1L4_8_Sn2L4_4,Sn1L4_9_Sn2L4_4,Sn1L4_10_Sn2L4_4,Sn1L4_11_Sn2L4_4,Sn1L4_12_Sn2L4_4,Sn1L4_13_Sn2L4_4,Sn1L4_14_Sn2L4_4,Sn1L4_15_Sn2L4_4,Sn1L4_16_Sn2L4_4,Sn1L4_17_Sn2L4_4,Sn1L4_18_Sn2L4_4,Sn1L4_19_Sn2L4_4,Sn1L4_20_Sn2L4_4,Sn1L4_21_Sn2L4_4,Sn1L4_22_Sn2L4_4,Sn1L4_23_Sn2L4_4,Sn1L4_24_Sn2L4_4,Sn1L4_25_Sn2L4_4,Sn1L4_26_Sn2L4_4,Sn1L4_27_Sn2L4_4,Sn1L4_28_Sn2L4_4: std_logic;
signal Sn1L5_4_Sn2L5_1,Sn1L5_5_Sn2L5_1,Sn1L5_6_Sn2L5_1,Sn1L5_7_Sn2L5_1,Sn1L5_8_Sn2L5_1,Sn1L5_9_Sn2L5_1,Sn1L5_10_Sn2L5_1,Sn1L5_11_Sn2L5_1,Sn1L5_12_Sn2L5_1,Sn1L5_13_Sn2L5_1,Sn1L5_14_Sn2L5_1,Sn1L5_15_Sn2L5_1,Sn1L5_16_Sn2L5_1,Sn1L5_17_Sn2L5_1,Sn1L5_18_Sn2L5_1,Sn1L5_19_Sn2L5_1,Sn1L5_20_Sn2L5_1,Sn1L5_21_Sn2L5_1,Sn1L5_22_Sn2L5_1,Sn1L5_23_Sn2L5_1,Sn1L5_24_Sn2L5_1,Sn1L5_25_Sn2L5_1,Sn1L5_26_Sn2L5_1,Sn1L5_27_Sn2L5_1,Sn1L5_28_Sn2L5_1,Sn1L5_29_Sn2L5_1:std_logic;
signal Sn1L5_5_Sn2L5_2,Sn1L5_6_Sn2L5_2,Sn1L5_7_Sn2L5_2,Sn1L5_8_Sn2L5_2,Sn1L5_9_Sn2L5_2,Sn1L5_10_Sn2L5_2,Sn1L5_11_Sn2L5_2,Sn1L5_12_Sn2L5_2,Sn1L5_13_Sn2L5_2,Sn1L5_14_Sn2L5_2,Sn1L5_15_Sn2L5_2,Sn1L5_16_Sn2L5_2,Sn1L5_17_Sn2L5_2,Sn1L5_18_Sn2L5_2,Sn1L5_19_Sn2L5_2,Sn1L5_20_Sn2L5_2,Sn1L5_21_Sn2L5_2,Sn1L5_22_Sn2L5_2,Sn1L5_23_Sn2L5_2,Sn1L5_24_Sn2L5_2,Sn1L5_25_Sn2L5_2,Sn1L5_26_Sn2L5_2,Sn1L5_27_Sn2L5_2,Sn1L5_28_Sn2L5_2,Sn1L5_29_Sn2L5_2,Sn1L5_30_Sn2L5_2:std_logic;
signal Sn1L6_3_Sn2L6_1,Sn1L6_4_Sn2L6_1,Sn1L6_5_Sn2L6_1,Sn1L6_6_Sn2L6_1,Sn1L6_7_Sn2L6_1,Sn1L6_8_Sn2L6_1,Sn1L6_9_Sn2L6_1,Sn1L6_10_Sn2L6_1,Sn1L6_11_Sn2L6_1,Sn1L6_12_Sn2L6_1,Sn1L6_13_Sn2L6_1,Sn1L6_14_Sn2L6_1,Sn1L6_15_Sn2L6_1,Sn1L6_16_Sn2L6_1,Sn1L6_17_Sn2L6_1,Sn1L6_18_Sn2L6_1,Sn1L6_19_Sn2L6_1,Sn1L6_20_Sn2L6_1,Sn1L6_21_Sn2L6_1,Sn1L6_22_Sn2L6_1,Sn1L6_23_Sn2L6_1,Sn1L6_24_Sn2L6_1,Sn1L6_25_Sn2L6_1,Sn1L6_26_Sn2L6_1,Sn1L6_27_Sn2L6_1,Sn1L6_28_Sn2L6_1,Sn1L6_29_Sn2L6_1,Sn1L6_30_Sn2L6_1:std_logic;
signal Sn1L6_4_Sn2L6_2,Sn1L6_5_Sn2L6_2,Sn1L6_6_Sn2L6_2,Sn1L6_7_Sn2L6_2,Sn1L6_8_Sn2L6_2,Sn1L6_9_Sn2L6_2,Sn1L6_10_Sn2L6_2,Sn1L6_11_Sn2L6_2,Sn1L6_12_Sn2L6_2,Sn1L6_13_Sn2L6_2,Sn1L6_14_Sn2L6_2,Sn1L6_15_Sn2L6_2,Sn1L6_16_Sn2L6_2,Sn1L6_17_Sn2L6_2,Sn1L6_18_Sn2L6_2,Sn1L6_19_Sn2L6_2,Sn1L6_20_Sn2L6_2,Sn1L6_21_Sn2L6_2,Sn1L6_22_Sn2L6_2,Sn1L6_23_Sn2L6_2,Sn1L6_24_Sn2L6_2,Sn1L6_25_Sn2L6_2,Sn1L6_26_Sn2L6_2,Sn1L6_27_Sn2L6_2,Sn1L6_28_Sn2L6_2,Sn1L6_29_Sn2L6_2,Sn1L6_30_Sn2L6_2,Sn1L6_31_Sn2L6_2:std_logic;

begin

dum0 <= A(0) nand B(0) after 150 ps;
A0B0 <= not dum0 after 100 ps;
dum1 <= A(0) nand B(1) after 150 ps;
A0B1 <= not dum1 after 100 ps;
dum2 <= A(1) nand B(0) after 150 ps;
A1B0 <= not dum2 after 100 ps;
dum3 <= A(0) nand B(2) after 150 ps;
A0B2 <= not dum3 after 100 ps;
dum4 <= A(1) nand B(1) after 150 ps;
A1B1 <= not dum4 after 100 ps;
dum5 <= A(2) nand B(0) after 150 ps;
A2B0 <= not dum5 after 100 ps;
dum6 <= A(0) nand B(3) after 150 ps;
A0B3 <= not dum6 after 100 ps;
dum7 <= A(1) nand B(2) after 150 ps;
A1B2 <= not dum7 after 100 ps;
dum8 <= A(2) nand B(1) after 150 ps;
A2B1 <= not dum8 after 100 ps;
dum9 <= A(3) nand B(0) after 150 ps;
A3B0 <= not dum9 after 100 ps;
dum10 <= A(0) nand B(4) after 150 ps;
A0B4 <= not dum10 after 100 ps;
dum11 <= A(1) nand B(3) after 150 ps;
A1B3 <= not dum11 after 100 ps;
dum12 <= A(2) nand B(2) after 150 ps;
A2B2 <= not dum12 after 100 ps;
dum13 <= A(3) nand B(1) after 150 ps;
A3B1 <= not dum13 after 100 ps;
dum14 <= A(4) nand B(0) after 150 ps;
A4B0 <= not dum14 after 100 ps;
dum15 <= A(0) nand B(5) after 150 ps;
A0B5 <= not dum15 after 100 ps;
dum16 <= A(1) nand B(4) after 150 ps;
A1B4 <= not dum16 after 100 ps;
dum17 <= A(2) nand B(3) after 150 ps;
A2B3 <= not dum17 after 100 ps;
dum18 <= A(3) nand B(2) after 150 ps;
A3B2 <= not dum18 after 100 ps;
dum19 <= A(4) nand B(1) after 150 ps;
A4B1 <= not dum19 after 100 ps;
dum20 <= A(5) nand B(0) after 150 ps;
A5B0 <= not dum20 after 100 ps;
dum21 <= A(0) nand B(6) after 150 ps;
A0B6 <= not dum21 after 100 ps;
dum22 <= A(1) nand B(5) after 150 ps;
A1B5 <= not dum22 after 100 ps;
dum23 <= A(2) nand B(4) after 150 ps;
A2B4 <= not dum23 after 100 ps;
dum24 <= A(3) nand B(3) after 150 ps;
A3B3 <= not dum24 after 100 ps;
dum25 <= A(4) nand B(2) after 150 ps;
A4B2 <= not dum25 after 100 ps;
dum26 <= A(5) nand B(1) after 150 ps;
A5B1 <= not dum26 after 100 ps;
dum27 <= A(6) nand B(0) after 150 ps;
A6B0 <= not dum27 after 100 ps;
dum28 <= A(0) nand B(7) after 150 ps;
A0B7 <= not dum28 after 100 ps;
dum29 <= A(1) nand B(6) after 150 ps;
A1B6 <= not dum29 after 100 ps;
dum30 <= A(2) nand B(5) after 150 ps;
A2B5 <= not dum30 after 100 ps;
dum31 <= A(3) nand B(4) after 150 ps;
A3B4 <= not dum31 after 100 ps;
dum32 <= A(4) nand B(3) after 150 ps;
A4B3 <= not dum32 after 100 ps;
dum33 <= A(5) nand B(2) after 150 ps;
A5B2 <= not dum33 after 100 ps;
dum34 <= A(6) nand B(1) after 150 ps;
A6B1 <= not dum34 after 100 ps;
dum35 <= A(7) nand B(0) after 150 ps;
A7B0 <= not dum35 after 100 ps;
dum36 <= A(0) nand B(8) after 150 ps;
A0B8 <= not dum36 after 100 ps;
dum37 <= A(1) nand B(7) after 150 ps;
A1B7 <= not dum37 after 100 ps;
dum38 <= A(2) nand B(6) after 150 ps;
A2B6 <= not dum38 after 100 ps;
dum39 <= A(3) nand B(5) after 150 ps;
A3B5 <= not dum39 after 100 ps;
dum40 <= A(4) nand B(4) after 150 ps;
A4B4 <= not dum40 after 100 ps;
dum41 <= A(5) nand B(3) after 150 ps;
A5B3 <= not dum41 after 100 ps;
dum42 <= A(6) nand B(2) after 150 ps;
A6B2 <= not dum42 after 100 ps;
dum43 <= A(7) nand B(1) after 150 ps;
A7B1 <= not dum43 after 100 ps;
dum44 <= A(8) nand B(0) after 150 ps;
A8B0 <= not dum44 after 100 ps;
dum45 <= A(0) nand B(9) after 150 ps;
A0B9 <= not dum45 after 100 ps;
dum46 <= A(1) nand B(8) after 150 ps;
A1B8 <= not dum46 after 100 ps;
dum47 <= A(2) nand B(7) after 150 ps;
A2B7 <= not dum47 after 100 ps;
dum48 <= A(3) nand B(6) after 150 ps;
A3B6 <= not dum48 after 100 ps;
dum49 <= A(4) nand B(5) after 150 ps;
A4B5 <= not dum49 after 100 ps;
dum50 <= A(5) nand B(4) after 150 ps;
A5B4 <= not dum50 after 100 ps;
dum51 <= A(6) nand B(3) after 150 ps;
A6B3 <= not dum51 after 100 ps;
dum52 <= A(7) nand B(2) after 150 ps;
A7B2 <= not dum52 after 100 ps;
dum53 <= A(8) nand B(1) after 150 ps;
A8B1 <= not dum53 after 100 ps;
dum54 <= A(9) nand B(0) after 150 ps;
A9B0 <= not dum54 after 100 ps;
dum55 <= A(0) nand B(10) after 150 ps;
A0B10 <= not dum55 after 100 ps;
dum56 <= A(1) nand B(9) after 150 ps;
A1B9 <= not dum56 after 100 ps;
dum57 <= A(2) nand B(8) after 150 ps;
A2B8 <= not dum57 after 100 ps;
dum58 <= A(3) nand B(7) after 150 ps;
A3B7 <= not dum58 after 100 ps;
dum59 <= A(4) nand B(6) after 150 ps;
A4B6 <= not dum59 after 100 ps;
dum60 <= A(5) nand B(5) after 150 ps;
A5B5 <= not dum60 after 100 ps;
dum61 <= A(6) nand B(4) after 150 ps;
A6B4 <= not dum61 after 100 ps;
dum62 <= A(7) nand B(3) after 150 ps;
A7B3 <= not dum62 after 100 ps;
dum63 <= A(8) nand B(2) after 150 ps;
A8B2 <= not dum63 after 100 ps;
dum64 <= A(9) nand B(1) after 150 ps;
A9B1 <= not dum64 after 100 ps;
dum65 <= A(10) nand B(0) after 150 ps;
A10B0 <= not dum65 after 100 ps;
dum66 <= A(0) nand B(11) after 150 ps;
A0B11 <= not dum66 after 100 ps;
dum67 <= A(1) nand B(10) after 150 ps;
A1B10 <= not dum67 after 100 ps;
dum68 <= A(2) nand B(9) after 150 ps;
A2B9 <= not dum68 after 100 ps;
dum69 <= A(3) nand B(8) after 150 ps;
A3B8 <= not dum69 after 100 ps;
dum70 <= A(4) nand B(7) after 150 ps;
A4B7 <= not dum70 after 100 ps;
dum71 <= A(5) nand B(6) after 150 ps;
A5B6 <= not dum71 after 100 ps;
dum72 <= A(6) nand B(5) after 150 ps;
A6B5 <= not dum72 after 100 ps;
dum73 <= A(7) nand B(4) after 150 ps;
A7B4 <= not dum73 after 100 ps;
dum74 <= A(8) nand B(3) after 150 ps;
A8B3 <= not dum74 after 100 ps;
dum75 <= A(9) nand B(2) after 150 ps;
A9B2 <= not dum75 after 100 ps;
dum76 <= A(10) nand B(1) after 150 ps;
A10B1 <= not dum76 after 100 ps;
dum77 <= A(11) nand B(0) after 150 ps;
A11B0 <= not dum77 after 100 ps;
dum78 <= A(0) nand B(12) after 150 ps;
A0B12 <= not dum78 after 100 ps;
dum79 <= A(1) nand B(11) after 150 ps;
A1B11 <= not dum79 after 100 ps;
dum80 <= A(2) nand B(10) after 150 ps;
A2B10 <= not dum80 after 100 ps;
dum81 <= A(3) nand B(9) after 150 ps;
A3B9 <= not dum81 after 100 ps;
dum82 <= A(4) nand B(8) after 150 ps;
A4B8 <= not dum82 after 100 ps;
dum83 <= A(5) nand B(7) after 150 ps;
A5B7 <= not dum83 after 100 ps;
dum84 <= A(6) nand B(6) after 150 ps;
A6B6 <= not dum84 after 100 ps;
dum85 <= A(7) nand B(5) after 150 ps;
A7B5 <= not dum85 after 100 ps;
dum86 <= A(8) nand B(4) after 150 ps;
A8B4 <= not dum86 after 100 ps;
dum87 <= A(9) nand B(3) after 150 ps;
A9B3 <= not dum87 after 100 ps;
dum88 <= A(10) nand B(2) after 150 ps;
A10B2 <= not dum88 after 100 ps;
dum89 <= A(11) nand B(1) after 150 ps;
A11B1 <= not dum89 after 100 ps;
dum90 <= A(12) nand B(0) after 150 ps;
A12B0 <= not dum90 after 100 ps;
dum91 <= A(0) nand B(13) after 150 ps;
A0B13 <= not dum91 after 100 ps;
dum92 <= A(1) nand B(12) after 150 ps;
A1B12 <= not dum92 after 100 ps;
dum93 <= A(2) nand B(11) after 150 ps;
A2B11 <= not dum93 after 100 ps;
dum94 <= A(3) nand B(10) after 150 ps;
A3B10 <= not dum94 after 100 ps;
dum95 <= A(4) nand B(9) after 150 ps;
A4B9 <= not dum95 after 100 ps;
dum96 <= A(5) nand B(8) after 150 ps;
A5B8 <= not dum96 after 100 ps;
dum97 <= A(6) nand B(7) after 150 ps;
A6B7 <= not dum97 after 100 ps;
dum98 <= A(7) nand B(6) after 150 ps;
A7B6 <= not dum98 after 100 ps;
dum99 <= A(8) nand B(5) after 150 ps;
A8B5 <= not dum99 after 100 ps;
dum100 <= A(9) nand B(4) after 150 ps;
A9B4 <= not dum100 after 100 ps;
dum101 <= A(10) nand B(3) after 150 ps;
A10B3 <= not dum101 after 100 ps;
dum102 <= A(11) nand B(2) after 150 ps;
A11B2 <= not dum102 after 100 ps;
dum103 <= A(12) nand B(1) after 150 ps;
A12B1 <= not dum103 after 100 ps;
dum104 <= A(13) nand B(0) after 150 ps;
A13B0 <= not dum104 after 100 ps;
dum105 <= A(0) nand B(14) after 150 ps;
A0B14 <= not dum105 after 100 ps;
dum106 <= A(1) nand B(13) after 150 ps;
A1B13 <= not dum106 after 100 ps;
dum107 <= A(2) nand B(12) after 150 ps;
A2B12 <= not dum107 after 100 ps;
dum108 <= A(3) nand B(11) after 150 ps;
A3B11 <= not dum108 after 100 ps;
dum109 <= A(4) nand B(10) after 150 ps;
A4B10 <= not dum109 after 100 ps;
dum110 <= A(5) nand B(9) after 150 ps;
A5B9 <= not dum110 after 100 ps;
dum111 <= A(6) nand B(8) after 150 ps;
A6B8 <= not dum111 after 100 ps;
dum112 <= A(7) nand B(7) after 150 ps;
A7B7 <= not dum112 after 100 ps;
dum113 <= A(8) nand B(6) after 150 ps;
A8B6 <= not dum113 after 100 ps;
dum114 <= A(9) nand B(5) after 150 ps;
A9B5 <= not dum114 after 100 ps;
dum115 <= A(10) nand B(4) after 150 ps;
A10B4 <= not dum115 after 100 ps;
dum116 <= A(11) nand B(3) after 150 ps;
A11B3 <= not dum116 after 100 ps;
dum117 <= A(12) nand B(2) after 150 ps;
A12B2 <= not dum117 after 100 ps;
dum118 <= A(13) nand B(1) after 150 ps;
A13B1 <= not dum118 after 100 ps;
dum119 <= A(14) nand B(0) after 150 ps;
A14B0 <= not dum119 after 100 ps;
dum120 <= A(0) nand B(15) after 150 ps;
A0B15 <= not dum120 after 100 ps;
dum121 <= A(1) nand B(14) after 150 ps;
A1B14 <= not dum121 after 100 ps;
dum122 <= A(2) nand B(13) after 150 ps;
A2B13 <= not dum122 after 100 ps;
dum123 <= A(3) nand B(12) after 150 ps;
A3B12 <= not dum123 after 100 ps;
dum124 <= A(4) nand B(11) after 150 ps;
A4B11 <= not dum124 after 100 ps;
dum125 <= A(5) nand B(10) after 150 ps;
A5B10 <= not dum125 after 100 ps;
dum126 <= A(6) nand B(9) after 150 ps;
A6B9 <= not dum126 after 100 ps;
dum127 <= A(7) nand B(8) after 150 ps;
A7B8 <= not dum127 after 100 ps;
dum128 <= A(8) nand B(7) after 150 ps;
A8B7 <= not dum128 after 100 ps;
dum129 <= A(9) nand B(6) after 150 ps;
A9B6 <= not dum129 after 100 ps;
dum130 <= A(10) nand B(5) after 150 ps;
A10B5 <= not dum130 after 100 ps;
dum131 <= A(11) nand B(4) after 150 ps;
A11B4 <= not dum131 after 100 ps;
dum132 <= A(12) nand B(3) after 150 ps;
A12B3 <= not dum132 after 100 ps;
dum133 <= A(13) nand B(2) after 150 ps;
A13B2 <= not dum133 after 100 ps;
dum134 <= A(14) nand B(1) after 150 ps;
A14B1 <= not dum134 after 100 ps;
dum135 <= A(15) nand B(0) after 150 ps;
A15B0 <= not dum135 after 100 ps;
dum136 <= A(1) nand B(15) after 150 ps;
A1B15 <= not dum136 after 100 ps;
dum137 <= A(2) nand B(14) after 150 ps;
A2B14 <= not dum137 after 100 ps;
dum138 <= A(3) nand B(13) after 150 ps;
A3B13 <= not dum138 after 100 ps;
dum139 <= A(4) nand B(12) after 150 ps;
A4B12 <= not dum139 after 100 ps;
dum140 <= A(5) nand B(11) after 150 ps;
A5B11 <= not dum140 after 100 ps;
dum141 <= A(6) nand B(10) after 150 ps;
A6B10 <= not dum141 after 100 ps;
dum142 <= A(7) nand B(9) after 150 ps;
A7B9 <= not dum142 after 100 ps;
dum143 <= A(8) nand B(8) after 150 ps;
A8B8 <= not dum143 after 100 ps;
dum144 <= A(9) nand B(7) after 150 ps;
A9B7 <= not dum144 after 100 ps;
dum145 <= A(10) nand B(6) after 150 ps;
A10B6 <= not dum145 after 100 ps;
dum146 <= A(11) nand B(5) after 150 ps;
A11B5 <= not dum146 after 100 ps;
dum147 <= A(12) nand B(4) after 150 ps;
A12B4 <= not dum147 after 100 ps;
dum148 <= A(13) nand B(3) after 150 ps;
A13B3 <= not dum148 after 100 ps;
dum149 <= A(14) nand B(2) after 150 ps;
A14B2 <= not dum149 after 100 ps;
dum150 <= A(15) nand B(1) after 150 ps;
A15B1 <= not dum150 after 100 ps;
dum151 <= A(2) nand B(15) after 150 ps;
A2B15 <= not dum151 after 100 ps;
dum152 <= A(3) nand B(14) after 150 ps;
A3B14 <= not dum152 after 100 ps;
dum153 <= A(4) nand B(13) after 150 ps;
A4B13 <= not dum153 after 100 ps;
dum154 <= A(5) nand B(12) after 150 ps;
A5B12 <= not dum154 after 100 ps;
dum155 <= A(6) nand B(11) after 150 ps;
A6B11 <= not dum155 after 100 ps;
dum156 <= A(7) nand B(10) after 150 ps;
A7B10 <= not dum156 after 100 ps;
dum157 <= A(8) nand B(9) after 150 ps;
A8B9 <= not dum157 after 100 ps;
dum158 <= A(9) nand B(8) after 150 ps;
A9B8 <= not dum158 after 100 ps;
dum159 <= A(10) nand B(7) after 150 ps;
A10B7 <= not dum159 after 100 ps;
dum160 <= A(11) nand B(6) after 150 ps;
A11B6 <= not dum160 after 100 ps;
dum161 <= A(12) nand B(5) after 150 ps;
A12B5 <= not dum161 after 100 ps;
dum162 <= A(13) nand B(4) after 150 ps;
A13B4 <= not dum162 after 100 ps;
dum163 <= A(14) nand B(3) after 150 ps;
A14B3 <= not dum163 after 100 ps;
dum164 <= A(15) nand B(2) after 150 ps;
A15B2 <= not dum164 after 100 ps;
dum165 <= A(3) nand B(15) after 150 ps;
A3B15 <= not dum165 after 100 ps;
dum166 <= A(4) nand B(14) after 150 ps;
A4B14 <= not dum166 after 100 ps;
dum167 <= A(5) nand B(13) after 150 ps;
A5B13 <= not dum167 after 100 ps;
dum168 <= A(6) nand B(12) after 150 ps;
A6B12 <= not dum168 after 100 ps;
dum169 <= A(7) nand B(11) after 150 ps;
A7B11 <= not dum169 after 100 ps;
dum170 <= A(8) nand B(10) after 150 ps;
A8B10 <= not dum170 after 100 ps;
dum171 <= A(9) nand B(9) after 150 ps;
A9B9 <= not dum171 after 100 ps;
dum172 <= A(10) nand B(8) after 150 ps;
A10B8 <= not dum172 after 100 ps;
dum173 <= A(11) nand B(7) after 150 ps;
A11B7 <= not dum173 after 100 ps;
dum174 <= A(12) nand B(6) after 150 ps;
A12B6 <= not dum174 after 100 ps;
dum175 <= A(13) nand B(5) after 150 ps;
A13B5 <= not dum175 after 100 ps;
dum176 <= A(14) nand B(4) after 150 ps;
A14B4 <= not dum176 after 100 ps;
dum177 <= A(15) nand B(3) after 150 ps;
A15B3 <= not dum177 after 100 ps;
dum178 <= A(4) nand B(15) after 150 ps;
A4B15 <= not dum178 after 100 ps;
dum179 <= A(5) nand B(14) after 150 ps;
A5B14 <= not dum179 after 100 ps;
dum180 <= A(6) nand B(13) after 150 ps;
A6B13 <= not dum180 after 100 ps;
dum181 <= A(7) nand B(12) after 150 ps;
A7B12 <= not dum181 after 100 ps;
dum182 <= A(8) nand B(11) after 150 ps;
A8B11 <= not dum182 after 100 ps;
dum183 <= A(9) nand B(10) after 150 ps;
A9B10 <= not dum183 after 100 ps;
dum184 <= A(10) nand B(9) after 150 ps;
A10B9 <= not dum184 after 100 ps;
dum185 <= A(11) nand B(8) after 150 ps;
A11B8 <= not dum185 after 100 ps;
dum186 <= A(12) nand B(7) after 150 ps;
A12B7 <= not dum186 after 100 ps;
dum187 <= A(13) nand B(6) after 150 ps;
A13B6 <= not dum187 after 100 ps;
dum188 <= A(14) nand B(5) after 150 ps;
A14B5 <= not dum188 after 100 ps;
dum189 <= A(15) nand B(4) after 150 ps;
A15B4 <= not dum189 after 100 ps;
dum190 <= A(5) nand B(15) after 150 ps;
A5B15 <= not dum190 after 100 ps;
dum191 <= A(6) nand B(14) after 150 ps;
A6B14 <= not dum191 after 100 ps;
dum192 <= A(7) nand B(13) after 150 ps;
A7B13 <= not dum192 after 100 ps;
dum193 <= A(8) nand B(12) after 150 ps;
A8B12 <= not dum193 after 100 ps;
dum194 <= A(9) nand B(11) after 150 ps;
A9B11 <= not dum194 after 100 ps;
dum195 <= A(10) nand B(10) after 150 ps;
A10B10 <= not dum195 after 100 ps;
dum196 <= A(11) nand B(9) after 150 ps;
A11B9 <= not dum196 after 100 ps;
dum197 <= A(12) nand B(8) after 150 ps;
A12B8 <= not dum197 after 100 ps;
dum198 <= A(13) nand B(7) after 150 ps;
A13B7 <= not dum198 after 100 ps;
dum199 <= A(14) nand B(6) after 150 ps;
A14B6 <= not dum199 after 100 ps;
dum200 <= A(15) nand B(5) after 150 ps;
A15B5 <= not dum200 after 100 ps;
dum201 <= A(6) nand B(15) after 150 ps;
A6B15 <= not dum201 after 100 ps;
dum202 <= A(7) nand B(14) after 150 ps;
A7B14 <= not dum202 after 100 ps;
dum203 <= A(8) nand B(13) after 150 ps;
A8B13 <= not dum203 after 100 ps;
dum204 <= A(9) nand B(12) after 150 ps;
A9B12 <= not dum204 after 100 ps;
dum205 <= A(10) nand B(11) after 150 ps;
A10B11 <= not dum205 after 100 ps;
dum206 <= A(11) nand B(10) after 150 ps;
A11B10 <= not dum206 after 100 ps;
dum207 <= A(12) nand B(9) after 150 ps;
A12B9 <= not dum207 after 100 ps;
dum208 <= A(13) nand B(8) after 150 ps;
A13B8 <= not dum208 after 100 ps;
dum209 <= A(14) nand B(7) after 150 ps;
A14B7 <= not dum209 after 100 ps;
dum210 <= A(15) nand B(6) after 150 ps;
A15B6 <= not dum210 after 100 ps;
dum211 <= A(7) nand B(15) after 150 ps;
A7B15 <= not dum211 after 100 ps;
dum212 <= A(8) nand B(14) after 150 ps;
A8B14 <= not dum212 after 100 ps;
dum213 <= A(9) nand B(13) after 150 ps;
A9B13 <= not dum213 after 100 ps;
dum214 <= A(10) nand B(12) after 150 ps;
A10B12 <= not dum214 after 100 ps;
dum215 <= A(11) nand B(11) after 150 ps;
A11B11 <= not dum215 after 100 ps;
dum216 <= A(12) nand B(10) after 150 ps;
A12B10 <= not dum216 after 100 ps;
dum217 <= A(13) nand B(9) after 150 ps;
A13B9 <= not dum217 after 100 ps;
dum218 <= A(14) nand B(8) after 150 ps;
A14B8 <= not dum218 after 100 ps;
dum219 <= A(15) nand B(7) after 150 ps;
A15B7 <= not dum219 after 100 ps;
dum220 <= A(8) nand B(15) after 150 ps;
A8B15 <= not dum220 after 100 ps;
dum221 <= A(9) nand B(14) after 150 ps;
A9B14 <= not dum221 after 100 ps;
dum222 <= A(10) nand B(13) after 150 ps;
A10B13 <= not dum222 after 100 ps;
dum223 <= A(11) nand B(12) after 150 ps;
A11B12 <= not dum223 after 100 ps;
dum224 <= A(12) nand B(11) after 150 ps;
A12B11 <= not dum224 after 100 ps;
dum225 <= A(13) nand B(10) after 150 ps;
A13B10 <= not dum225 after 100 ps;
dum226 <= A(14) nand B(9) after 150 ps;
A14B9 <= not dum226 after 100 ps;
dum227 <= A(15) nand B(8) after 150 ps;
A15B8 <= not dum227 after 100 ps;
dum228 <= A(9) nand B(15) after 150 ps;
A9B15 <= not dum228 after 100 ps;
dum229 <= A(10) nand B(14) after 150 ps;
A10B14 <= not dum229 after 100 ps;
dum230 <= A(11) nand B(13) after 150 ps;
A11B13 <= not dum230 after 100 ps;
dum231 <= A(12) nand B(12) after 150 ps;
A12B12 <= not dum231 after 100 ps;
dum232 <= A(13) nand B(11) after 150 ps;
A13B11 <= not dum232 after 100 ps;
dum233 <= A(14) nand B(10) after 150 ps;
A14B10 <= not dum233 after 100 ps;
dum234 <= A(15) nand B(9) after 150 ps;
A15B9 <= not dum234 after 100 ps;
dum235 <= A(10) nand B(15) after 150 ps;
A10B15 <= not dum235 after 100 ps;
dum236 <= A(11) nand B(14) after 150 ps;
A11B14 <= not dum236 after 100 ps;
dum237 <= A(12) nand B(13) after 150 ps;
A12B13 <= not dum237 after 100 ps;
dum238 <= A(13) nand B(12) after 150 ps;
A13B12 <= not dum238 after 100 ps;
dum239 <= A(14) nand B(11) after 150 ps;
A14B11 <= not dum239 after 100 ps;
dum240 <= A(15) nand B(10) after 150 ps;
A15B10 <= not dum240 after 100 ps;
dum241 <= A(11) nand B(15) after 150 ps;
A11B15 <= not dum241 after 100 ps;
dum242 <= A(12) nand B(14) after 150 ps;
A12B14 <= not dum242 after 100 ps;
dum243 <= A(13) nand B(13) after 150 ps;
A13B13 <= not dum243 after 100 ps;
dum244 <= A(14) nand B(12) after 150 ps;
A14B12 <= not dum244 after 100 ps;
dum245 <= A(15) nand B(11) after 150 ps;
A15B11 <= not dum245 after 100 ps;
dum246 <= A(12) nand B(15) after 150 ps;
A12B15 <= not dum246 after 100 ps;
dum247 <= A(13) nand B(14) after 150 ps;
A13B14 <= not dum247 after 100 ps;
dum248 <= A(14) nand B(13) after 150 ps;
A14B13 <= not dum248 after 100 ps;
dum249 <= A(15) nand B(12) after 150 ps;
A15B12 <= not dum249 after 100 ps;
dum250 <= A(13) nand B(15) after 150 ps;
A13B15 <= not dum250 after 100 ps;
dum251 <= A(14) nand B(14) after 150 ps;
A14B14 <= not dum251 after 100 ps;
dum252 <= A(15) nand B(13) after 150 ps;
A15B13 <= not dum252 after 100 ps;
dum253 <= A(14) nand B(15) after 150 ps;
A14B15 <= not dum253 after 100 ps;
dum254 <= A(15) nand B(14) after 150 ps;
A15B14 <= not dum254 after 100 ps;
dum255 <= A(15) nand B(15) after 150 ps;
A15B15 <= not dum255 after 100 ps;

HALFADD_01: HALFADD port map (A13B0,A12B1,Sn1L1_14_Sn2L1_1,Sn1L1_15_Sn2L1_2);
HALFADD_02: HALFADD port map (A14B0,A13B1,Sn1L1_15_Sn2L1_1,Sn1L1_16_Sn2L1_2);
HALFADD_03: HALFADD port map (A15B0,A14B1,Sn1L1_16_Sn2L1_1,Sn1L1_17_Sn2L1_2);
HALFADD_04: HALFADD port map (A15B1,A14B2,Sn1L1_17_Sn2L1_1,Sn1L1_18_Sn2L1_2);

FULLADD_01: FULLADD port map (A12B2,A11B3,A10B4,Sn1L1_15_Sn2L1_3,Sn1L1_16_Sn2L1_4);
FULLADD_02: FULLADD port map (A13B2,A12B3,A11B4,Sn1L1_16_Sn2L1_3,Sn1L1_17_Sn2L1_4);
FULLADD_03: FULLADD port map (A10B5,A9B6,A8B7,Sn1L1_16_Sn2L1_5,Sn1L1_17_Sn2L1_6);
FULLADD_04: FULLADD port map (A13B3,A12B4,A11B5,Sn1L1_17_Sn2L1_3,Sn1L1_18_Sn2L1_4);
FULLADD_05: FULLADD port map (A10B6,A9B7,A8B8,Sn1L1_17_Sn2L1_5,Sn1L1_18_Sn2L1_6);
FULLADD_06: FULLADD port map (A15B2,A14B3,A13B4,Sn1L1_18_Sn2L1_1,Sn1L1_19_Sn2L1_2);
FULLADD_07: FULLADD port map (A12B5,A11B6,A10B7,Sn1L1_18_Sn2L1_3,Sn1L1_19_Sn2L1_4);
FULLADD_08: FULLADD port map (A15B3,A14B4,A13B5,Sn1L1_19_Sn2L1_1,Sn1L1_20_Sn2L1_2);

HALFADD_05: HALFADD port map (A9B0,A8B1,Sn1L2_10_Sn2L2_1,Sn1L2_11_Sn2L2_2);
HALFADD_06: HALFADD port map (A10B0,A9B1,Sn1L2_11_Sn2L2_1,Sn1L2_12_Sn2L2_2);
HALFADD_07: HALFADD port map (A11B0,A10B1,Sn1L2_12_Sn2L2_1,Sn1L2_13_Sn2L2_2);
HALFADD_08: HALFADD port map (A12B0,A11B1,Sn1L2_13_Sn2L2_1,Sn1L2_14_Sn2L2_2);
FULLADD_09: FULLADD port map (A8B2,A7B3,A6B4,Sn1L2_11_Sn2L2_3,Sn1L2_12_Sn2L2_4);
FULLADD_10: FULLADD port map (A9B2,A8B3,A7B4,Sn1L2_12_Sn2L2_3,Sn1L2_13_Sn2L2_4);
FULLADD_11: FULLADD port map (A6B5,A5B6,A4B7,Sn1L2_12_Sn2L2_5,Sn1L2_13_Sn2L2_6);
FULLADD_12: FULLADD port map (A10B2,A9B3,A8B4,Sn1L2_13_Sn2L2_3,Sn1L2_14_Sn2L2_4);
FULLADD_13: FULLADD port map (A7B5,A6B6,A5B7,Sn1L2_13_Sn2L2_5,Sn1L2_14_Sn2L2_6);
FULLADD_14: FULLADD port map (A4B8,A3B9,A2B10,Sn1L2_13_Sn2L2_7,Sn1L2_14_Sn2L2_8);
FULLADD_15: FULLADD port map (Sn1L1_14_Sn2L1_1,A11B2,A10B3,Sn1L2_14_Sn2L2_1,Sn1L2_15_Sn2L2_2);
FULLADD_16: FULLADD port map (Sn1L1_15_Sn2L1_1,Sn1L1_15_Sn2L1_2,Sn1L1_15_Sn2L1_3,Sn1L2_15_Sn2L2_1,Sn1L2_16_Sn2L2_2);
FULLADD_17: FULLADD port map (Sn1L1_16_Sn2L1_1,Sn1L1_16_Sn2L1_2,Sn1L1_16_Sn2L1_3,Sn1L2_16_Sn2L2_1,Sn1L2_17_Sn2L2_2);
FULLADD_18: FULLADD port map (Sn1L1_17_Sn2L1_1,Sn1L1_17_Sn2L1_2,Sn1L1_17_Sn2L1_3,Sn1L2_17_Sn2L2_1,Sn1L2_18_Sn2L2_2);
FULLADD_19: FULLADD port map (Sn1L1_18_Sn2L1_1,Sn1L1_18_Sn2L1_2,Sn1L1_18_Sn2L1_3,Sn1L2_18_Sn2L2_1,Sn1L2_19_Sn2L2_2);
FULLADD_20: FULLADD port map (Sn1L1_19_Sn2L1_1,Sn1L1_19_Sn2L1_2,A12B6,Sn1L2_19_Sn2L2_1,Sn1L2_20_Sn2L2_2);
FULLADD_21: FULLADD port map (A15B4,Sn1L1_20_Sn2L1_2,A14B5,Sn1L2_20_Sn2L2_1,Sn1L2_21_Sn2L2_2);
FULLADD_22: FULLADD port map (A15B5,A14B6,A13B7,Sn1L2_21_Sn2L2_1,Sn1L2_22_Sn2L2_2);
FULLADD_23: FULLADD port map (A15B6,A14B7,A13B8,Sn1L2_22_Sn2L2_1,Sn1L2_23_Sn2L2_2);
FULLADD_24: FULLADD port map (A15B7,A14B8,A13B9,Sn1L2_23_Sn2L2_1,Sn1L2_24_Sn2L2_2);
FULLADD_25: FULLADD port map (A9B4,A8B5,A7B6,Sn1L2_14_Sn2L2_3,Sn1L2_15_Sn2L2_4);
FULLADD_26: FULLADD port map (A9B5,A8B6,A7B7,Sn1L2_15_Sn2L2_3,Sn1L2_16_Sn2L2_4);
FULLADD_27: FULLADD port map (Sn1L1_16_Sn2L1_4,Sn1L1_16_Sn2L1_5,A7B8,Sn1L2_16_Sn2L2_3,Sn1L2_17_Sn2L2_4);
FULLADD_28: FULLADD port map (Sn1L1_17_Sn2L1_4,Sn1L1_17_Sn2L1_5,Sn1L1_17_Sn2L1_6,Sn1L2_17_Sn2L2_3,Sn1L2_18_Sn2L2_4);
FULLADD_29: FULLADD port map (Sn1L1_18_Sn2L1_4,A9B8,Sn1L1_18_Sn2L1_6,Sn1L2_18_Sn2L2_3,Sn1L2_19_Sn2L2_4);
FULLADD_30: FULLADD port map (Sn1L1_19_Sn2L1_4,A11B7,A10B8,Sn1L2_19_Sn2L2_3,Sn1L2_20_Sn2L2_4);
FULLADD_31: FULLADD port map (A13B6,A12B7,A11B8,Sn1L2_20_Sn2L2_3,Sn1L2_21_Sn2L2_4);
FULLADD_32: FULLADD port map (A12B8,A11B9,A10B10,Sn1L2_21_Sn2L2_3,Sn1L2_22_Sn2L2_4);
FULLADD_33: FULLADD port map (A12B9,A11B10,A10B11,Sn1L2_22_Sn2L2_3,Sn1L2_23_Sn2L2_4);
FULLADD_34: FULLADD port map (A6B7,A5B8,A4B9,Sn1L2_14_Sn2L2_5,Sn1L2_15_Sn2L2_6);
FULLADD_35: FULLADD port map (A6B8,A5B9,A4B10,Sn1L2_15_Sn2L2_5,Sn1L2_16_Sn2L2_6);
FULLADD_36: FULLADD port map (A6B9,A5B10,A4B11,Sn1L2_16_Sn2L2_5,Sn1L2_17_Sn2L2_6);
FULLADD_37: FULLADD port map (A7B9,A6B10,A5B11,Sn1L2_17_Sn2L2_5,Sn1L2_18_Sn2L2_6);
FULLADD_38: FULLADD port map (A8B9,A7B10,A6B11,Sn1L2_18_Sn2L2_5,Sn1L2_19_Sn2L2_6);
FULLADD_39: FULLADD port map (A9B9,A8B10,A7B11,Sn1L2_19_Sn2L2_5,Sn1L2_20_Sn2L2_6);
FULLADD_40: FULLADD port map (A10B9,A9B10,A8B11,Sn1L2_20_Sn2L2_5,Sn1L2_21_Sn2L2_6);
FULLADD_41: FULLADD port map (A9B11,A8B12,A7B13,Sn1L2_21_Sn2L2_5,Sn1L2_22_Sn2L2_6);
FULLADD_42: FULLADD port map (A3B10,A2B11,A1B12,Sn1L2_14_Sn2L2_7,Sn1L2_15_Sn2L2_8);
FULLADD_43: FULLADD port map (A3B11,A2B12,A1B13,Sn1L2_15_Sn2L2_7,Sn1L2_16_Sn2L2_8);
FULLADD_44: FULLADD port map (A3B12,A2B13,A1B14,Sn1L2_16_Sn2L2_7,Sn1L2_17_Sn2L2_8);
FULLADD_45: FULLADD port map (A4B12,A3B13,A2B14,Sn1L2_17_Sn2L2_7,Sn1L2_18_Sn2L2_8);
FULLADD_46: FULLADD port map (A5B12,A4B13,A3B14,Sn1L2_18_Sn2L2_7,Sn1L2_19_Sn2L2_8);
FULLADD_47: FULLADD port map (A6B12,A5B13,A4B14,Sn1L2_19_Sn2L2_7,Sn1L2_20_Sn2L2_8);
FULLADD_48: FULLADD port map (A7B12,A6B13,A5B14,Sn1L2_20_Sn2L2_7,Sn1L2_21_Sn2L2_8);

HALFADD_9: HALFADD port map (A6B0,A5B1,Sn1L3_7_Sn2L3_1,Sn1L3_8_Sn2L3_2);
HALFADD_10: HALFADD port map (A7B0,A6B1,Sn1L3_8_Sn2L3_1,Sn1L3_9_Sn2L3_2);
HALFADD_11: HALFADD port map (A8B0,A7B1,Sn1L3_9_Sn2L3_1,Sn1L3_10_Sn2L3_2);

FULLADD_49: FULLADD port map (A5B2,A4B3,A3B4,Sn1L3_8_Sn2L3_3,Sn1L3_9_Sn2L3_4);
FULLADD_50: FULLADD port map (A6B2,A5B3,A4B4,Sn1L3_9_Sn2L3_3,Sn1L3_10_Sn2L3_4);
FULLADD_51: FULLADD port map (A3B5,A2B6,A1B7,Sn1L3_9_Sn2L3_5,Sn1L3_10_Sn2L3_6);
FULLADD_52: FULLADD port map (Sn1L2_10_Sn2L2_1,A7B2,A6B3,Sn1L3_10_Sn2L3_1,Sn1L3_11_Sn2L3_2);
FULLADD_53: FULLADD port map (Sn1L2_11_Sn2L2_1,Sn1L2_11_Sn2L2_2,Sn1L2_11_Sn2L2_3,Sn1L3_11_Sn2L3_1,Sn1L3_12_Sn2L3_2);
FULLADD_54: FULLADD port map (Sn1L2_12_Sn2L2_1,Sn1L2_12_Sn2L2_2,Sn1L2_12_Sn2L2_3,Sn1L3_12_Sn2L3_1,Sn1L3_13_Sn2L3_2);
FULLADD_55: FULLADD port map (Sn1L2_13_Sn2L2_1,Sn1L2_13_Sn2L2_2,Sn1L2_13_Sn2L2_3,Sn1L3_13_Sn2L3_1,Sn1L3_14_Sn2L3_2);
FULLADD_56: FULLADD port map (Sn1L2_14_Sn2L2_1,Sn1L2_14_Sn2L2_2,Sn1L2_14_Sn2L2_3,Sn1L3_14_Sn2L3_1,Sn1L3_15_Sn2L3_2);
FULLADD_57: FULLADD port map (Sn1L2_15_Sn2L2_1,Sn1L2_15_Sn2L2_2,Sn1L2_15_Sn2L2_3,Sn1L3_15_Sn2L3_1,Sn1L3_16_Sn2L3_2);
FULLADD_58: FULLADD port map (Sn1L2_16_Sn2L2_1,Sn1L2_16_Sn2L2_2,Sn1L2_16_Sn2L2_3,Sn1L3_16_Sn2L3_1,Sn1L3_17_Sn2L3_2);
FULLADD_59: FULLADD port map (Sn1L2_17_Sn2L2_1,Sn1L2_17_Sn2L2_2,Sn1L2_17_Sn2L2_3,Sn1L3_17_Sn2L3_1,Sn1L3_18_Sn2L3_2);
FULLADD_60: FULLADD port map (Sn1L2_18_Sn2L2_1,Sn1L2_18_Sn2L2_2,Sn1L2_18_Sn2L2_3,Sn1L3_18_Sn2L3_1,Sn1L3_19_Sn2L3_2);
FULLADD_61: FULLADD port map (Sn1L2_19_Sn2L2_1,Sn1L2_19_Sn2L2_2,Sn1L2_19_Sn2L2_3,Sn1L3_19_Sn2L3_1,Sn1L3_20_Sn2L3_2);
FULLADD_62: FULLADD port map (Sn1L2_20_Sn2L2_1,Sn1L2_20_Sn2L2_2,Sn1L2_20_Sn2L2_3,Sn1L3_20_Sn2L3_1,Sn1L3_21_Sn2L3_2);
FULLADD_63: FULLADD port map (Sn1L2_21_Sn2L2_1,Sn1L2_21_Sn2L2_2,Sn1L2_21_Sn2L2_3,Sn1L3_21_Sn2L3_1,Sn1L3_22_Sn2L3_2);
FULLADD_64: FULLADD port map (Sn1L2_22_Sn2L2_1,Sn1L2_22_Sn2L2_2,Sn1L2_22_Sn2L2_3,Sn1L3_22_Sn2L3_1,Sn1L3_23_Sn2L3_2);
FULLADD_65: FULLADD port map (Sn1L2_23_Sn2L2_1,Sn1L2_23_Sn2L2_2,A12B10,Sn1L3_23_Sn2L3_1,Sn1L3_24_Sn2L3_2);
FULLADD_66: FULLADD port map (A15B8,Sn1L2_24_Sn2L2_2,A14B9,Sn1L3_24_Sn2L3_1,Sn1L3_25_Sn2L3_2);
FULLADD_67: FULLADD port map (A15B9,A14B10,A13B11,Sn1L3_25_Sn2L3_1,Sn1L3_26_Sn2L3_2);
FULLADD_68: FULLADD port map (A15B10,A14B11,A13B12,Sn1L3_26_Sn2L3_1,Sn1L3_27_Sn2L3_2);
FULLADD_69: FULLADD port map (A5B4,A4B5,A3B6,Sn1L3_10_Sn2L3_3,Sn1L3_11_Sn2L3_4);
FULLADD_70: FULLADD port map (A5B5,A4B6,A3B7,Sn1L3_11_Sn2L3_3,Sn1L3_12_Sn2L3_4);
FULLADD_71: FULLADD port map (Sn1L2_12_Sn2L2_4,Sn1L2_12_Sn2L2_5,A3B8,Sn1L3_12_Sn2L3_3,Sn1L3_13_Sn2L3_4);
FULLADD_72: FULLADD port map (Sn1L2_13_Sn2L2_4,Sn1L2_13_Sn2L2_5,Sn1L2_13_Sn2L2_6,Sn1L3_13_Sn2L3_3,Sn1L3_14_Sn2L3_4);
FULLADD_73: FULLADD port map (Sn1L2_14_Sn2L2_4,Sn1L2_14_Sn2L2_5,Sn1L2_14_Sn2L2_6,Sn1L3_14_Sn2L3_3,Sn1L3_15_Sn2L3_4);
FULLADD_74: FULLADD port map (Sn1L2_15_Sn2L2_4,Sn1L2_15_Sn2L2_5,Sn1L2_15_Sn2L2_6,Sn1L3_15_Sn2L3_3,Sn1L3_16_Sn2L3_4);
FULLADD_75: FULLADD port map (Sn1L2_16_Sn2L2_4,Sn1L2_16_Sn2L2_5,Sn1L2_16_Sn2L2_6,Sn1L3_16_Sn2L3_3,Sn1L3_17_Sn2L3_4);
FULLADD_76: FULLADD port map (Sn1L2_17_Sn2L2_4,Sn1L2_17_Sn2L2_5,Sn1L2_17_Sn2L2_6,Sn1L3_17_Sn2L3_3,Sn1L3_18_Sn2L3_4);
FULLADD_77: FULLADD port map (Sn1L2_18_Sn2L2_4,Sn1L2_18_Sn2L2_5,Sn1L2_18_Sn2L2_6,Sn1L3_18_Sn2L3_3,Sn1L3_19_Sn2L3_4);
FULLADD_78: FULLADD port map (Sn1L2_19_Sn2L2_4,Sn1L2_19_Sn2L2_5,Sn1L2_19_Sn2L2_6,Sn1L3_19_Sn2L3_3,Sn1L3_20_Sn2L3_4);
FULLADD_79: FULLADD port map (Sn1L2_20_Sn2L2_4,Sn1L2_20_Sn2L2_5,Sn1L2_20_Sn2L2_6,Sn1L3_20_Sn2L3_3,Sn1L3_21_Sn2L3_4);
FULLADD_80: FULLADD port map (Sn1L2_21_Sn2L2_4,Sn1L2_21_Sn2L2_5,Sn1L2_21_Sn2L2_6,Sn1L3_21_Sn2L3_3,Sn1L3_22_Sn2L3_4);
FULLADD_81: FULLADD port map (Sn1L2_22_Sn2L2_4,A9B12,Sn1L2_22_Sn2L2_6,Sn1L3_22_Sn2L3_3,Sn1L3_23_Sn2L3_4);
FULLADD_82: FULLADD port map (Sn1L2_23_Sn2L2_4,A11B11,A10B12,Sn1L3_23_Sn2L3_3,Sn1L3_24_Sn2L3_4);
FULLADD_83: FULLADD port map (A13B10,A12B11,A11B12,Sn1L3_24_Sn2L3_3,Sn1L3_25_Sn2L3_4);
FULLADD_84: FULLADD port map (A12B12,A11B13,A10B14,Sn1L3_25_Sn2L3_3,Sn1L3_26_Sn2L3_4);
FULLADD_85: FULLADD port map (A2B7,A1B8,A0B9,Sn1L3_10_Sn2L3_5,Sn1L3_11_Sn2L3_6);
FULLADD_86: FULLADD port map (A2B8,A1B9,A0B10,Sn1L3_11_Sn2L3_5,Sn1L3_12_Sn2L3_6);
FULLADD_87: FULLADD port map (A2B9,A1B10,A0B11,Sn1L3_12_Sn2L3_5,Sn1L3_13_Sn2L3_6);
FULLADD_88: FULLADD port map (Sn1L2_13_Sn2L2_7,A1B11,A0B12,Sn1L3_13_Sn2L3_5,Sn1L3_14_Sn2L3_6);
FULLADD_89: FULLADD port map (Sn1L2_14_Sn2L2_7,Sn1L2_14_Sn2L2_8,A0B13,Sn1L3_14_Sn2L3_5,Sn1L3_15_Sn2L3_6);
FULLADD_90: FULLADD port map (Sn1L2_15_Sn2L2_7,Sn1L2_15_Sn2L2_8,A0B14,Sn1L3_15_Sn2L3_5,Sn1L3_16_Sn2L3_6);
FULLADD_91: FULLADD port map (Sn1L2_16_Sn2L2_7,Sn1L2_16_Sn2L2_8,A0B15,Sn1L3_16_Sn2L3_5,Sn1L3_17_Sn2L3_6);
FULLADD_92: FULLADD port map (Sn1L2_17_Sn2L2_7,Sn1L2_17_Sn2L2_8,A1B15,Sn1L3_17_Sn2L3_5,Sn1L3_18_Sn2L3_6);
FULLADD_93: FULLADD port map (Sn1L2_18_Sn2L2_7,Sn1L2_18_Sn2L2_8,A2B15,Sn1L3_18_Sn2L3_5,Sn1L3_19_Sn2L3_6);
FULLADD_94: FULLADD port map (Sn1L2_19_Sn2L2_7,Sn1L2_19_Sn2L2_8,A3B15,Sn1L3_19_Sn2L3_5,Sn1L3_20_Sn2L3_6);
FULLADD_95: FULLADD port map (Sn1L2_20_Sn2L2_7,Sn1L2_20_Sn2L2_8,A4B15,Sn1L3_20_Sn2L3_5,Sn1L3_21_Sn2L3_6);
FULLADD_96: FULLADD port map (A6B14,Sn1L2_21_Sn2L2_8,A5B15,Sn1L3_21_Sn2L3_5,Sn1L3_22_Sn2L3_6);
FULLADD_97: FULLADD port map (A8B13,A7B14,A6B15,Sn1L3_22_Sn2L3_5,Sn1L3_23_Sn2L3_6);
FULLADD_98: FULLADD port map (A9B13,A8B14,A7B15,Sn1L3_23_Sn2L3_5,Sn1L3_24_Sn2L3_6);
FULLADD_99: FULLADD port map (A10B13,A9B14,A8B15,Sn1L3_24_Sn2L3_5,Sn1L3_25_Sn2L3_6);

HALFADD_12: HALFADD port map (A4B0,A3B1,Sn1L4_5_Sn2L4_1,Sn1L4_6_Sn2L4_2);
HALFADD_13: HALFADD port map (A5B0,A4B1,Sn1L4_6_Sn2L4_1,Sn1L4_7_Sn2L4_2);

FULLADD_100: FULLADD port map (A3B2,A2B3,A1B4,Sn1L4_6_Sn2L4_3,Sn1L4_7_Sn2L4_4);
FULLADD_101: FULLADD port map (Sn1L3_7_Sn2L3_1,A4B2,A3B3,Sn1L4_7_Sn2L4_1,Sn1L4_8_Sn2L4_2);
FULLADD_102: FULLADD port map (Sn1L3_8_Sn2L3_1,Sn1L3_8_Sn2L3_2,Sn1L3_8_Sn2L3_3,Sn1L4_8_Sn2L4_1,Sn1L4_9_Sn2L4_2);
FULLADD_103: FULLADD port map (Sn1L3_9_Sn2L3_1,Sn1L3_9_Sn2L3_2,Sn1L3_9_Sn2L3_3,Sn1L4_9_Sn2L4_1,Sn1L4_10_Sn2L4_2);
FULLADD_104: FULLADD port map (Sn1L3_10_Sn2L3_1,Sn1L3_10_Sn2L3_2,Sn1L3_10_Sn2L3_3,Sn1L4_10_Sn2L4_1,Sn1L4_11_Sn2L4_2);
FULLADD_105: FULLADD port map (Sn1L3_11_Sn2L3_1,Sn1L3_11_Sn2L3_2,Sn1L3_11_Sn2L3_3,Sn1L4_11_Sn2L4_1,Sn1L4_12_Sn2L4_2);
FULLADD_106: FULLADD port map (Sn1L3_12_Sn2L3_1,Sn1L3_12_Sn2L3_2,Sn1L3_12_Sn2L3_3,Sn1L4_12_Sn2L4_1,Sn1L4_13_Sn2L4_2);
FULLADD_107: FULLADD port map (Sn1L3_13_Sn2L3_1,Sn1L3_13_Sn2L3_2,Sn1L3_13_Sn2L3_3,Sn1L4_13_Sn2L4_1,Sn1L4_14_Sn2L4_2);
FULLADD_108: FULLADD port map (Sn1L3_14_Sn2L3_1,Sn1L3_14_Sn2L3_2,Sn1L3_14_Sn2L3_3,Sn1L4_14_Sn2L4_1,Sn1L4_15_Sn2L4_2);
FULLADD_109: FULLADD port map (Sn1L3_15_Sn2L3_1,Sn1L3_15_Sn2L3_2,Sn1L3_15_Sn2L3_3,Sn1L4_15_Sn2L4_1,Sn1L4_16_Sn2L4_2);
FULLADD_110: FULLADD port map (Sn1L3_16_Sn2L3_1,Sn1L3_16_Sn2L3_2,Sn1L3_16_Sn2L3_3,Sn1L4_16_Sn2L4_1,Sn1L4_17_Sn2L4_2);
FULLADD_111: FULLADD port map (Sn1L3_17_Sn2L3_1,Sn1L3_17_Sn2L3_2,Sn1L3_17_Sn2L3_3,Sn1L4_17_Sn2L4_1,Sn1L4_18_Sn2L4_2);
FULLADD_112: FULLADD port map (Sn1L3_18_Sn2L3_1,Sn1L3_18_Sn2L3_2,Sn1L3_18_Sn2L3_3,Sn1L4_18_Sn2L4_1,Sn1L4_19_Sn2L4_2);
FULLADD_113: FULLADD port map (Sn1L3_19_Sn2L3_1,Sn1L3_19_Sn2L3_2,Sn1L3_19_Sn2L3_3,Sn1L4_19_Sn2L4_1,Sn1L4_20_Sn2L4_2);
FULLADD_114: FULLADD port map (Sn1L3_20_Sn2L3_1,Sn1L3_20_Sn2L3_2,Sn1L3_20_Sn2L3_3,Sn1L4_20_Sn2L4_1,Sn1L4_21_Sn2L4_2);
FULLADD_115: FULLADD port map (Sn1L3_21_Sn2L3_1,Sn1L3_21_Sn2L3_2,Sn1L3_21_Sn2L3_3,Sn1L4_21_Sn2L4_1,Sn1L4_22_Sn2L4_2);
FULLADD_116: FULLADD port map (Sn1L3_22_Sn2L3_1,Sn1L3_22_Sn2L3_2,Sn1L3_22_Sn2L3_3,Sn1L4_22_Sn2L4_1,Sn1L4_23_Sn2L4_2);
FULLADD_117: FULLADD port map (Sn1L3_23_Sn2L3_1,Sn1L3_23_Sn2L3_2,Sn1L3_23_Sn2L3_3,Sn1L4_23_Sn2L4_1,Sn1L4_24_Sn2L4_2);
FULLADD_118: FULLADD port map (Sn1L3_24_Sn2L3_1,Sn1L3_24_Sn2L3_2,Sn1L3_24_Sn2L3_3,Sn1L4_24_Sn2L4_1,Sn1L4_25_Sn2L4_2);
FULLADD_119: FULLADD port map (Sn1L3_25_Sn2L3_1,Sn1L3_25_Sn2L3_2,Sn1L3_25_Sn2L3_3,Sn1L4_25_Sn2L4_1,Sn1L4_26_Sn2L4_2);
FULLADD_120: FULLADD port map (Sn1L3_26_Sn2L3_1,Sn1L3_26_Sn2L3_2,A12B13,Sn1L4_26_Sn2L4_1,Sn1L4_27_Sn2L4_2);
FULLADD_121: FULLADD port map (A15B11,Sn1L3_27_Sn2L3_2,A14B12,Sn1L4_27_Sn2L4_1,Sn1L4_28_Sn2L4_2);
FULLADD_122: FULLADD port map (A15B12,A14B13,A13B14,Sn1L4_28_Sn2L4_1,Sn1L4_29_Sn2L4_2);
FULLADD_123: FULLADD port map (A2B4,A1B5,A0B6,Sn1L4_7_Sn2L4_3,Sn1L4_8_Sn2L4_4);
FULLADD_124: FULLADD port map (A2B5,A1B6,A0B7,Sn1L4_8_Sn2L4_3,Sn1L4_9_Sn2L4_4);
FULLADD_125: FULLADD port map (Sn1L3_9_Sn2L3_4,Sn1L3_9_Sn2L3_5,A0B8,Sn1L4_9_Sn2L4_3,Sn1L4_10_Sn2L4_4);
FULLADD_126: FULLADD port map (Sn1L3_10_Sn2L3_4,Sn1L3_10_Sn2L3_5,Sn1L3_10_Sn2L3_6,Sn1L4_10_Sn2L4_3,Sn1L4_11_Sn2L4_4);
FULLADD_127: FULLADD port map (Sn1L3_11_Sn2L3_4,Sn1L3_11_Sn2L3_5,Sn1L3_11_Sn2L3_6,Sn1L4_11_Sn2L4_3,Sn1L4_12_Sn2L4_4);
FULLADD_128: FULLADD port map (Sn1L3_12_Sn2L3_4,Sn1L3_12_Sn2L3_5,Sn1L3_12_Sn2L3_6,Sn1L4_12_Sn2L4_3,Sn1L4_13_Sn2L4_4);
FULLADD_129: FULLADD port map (Sn1L3_13_Sn2L3_4,Sn1L3_13_Sn2L3_5,Sn1L3_13_Sn2L3_6,Sn1L4_13_Sn2L4_3,Sn1L4_14_Sn2L4_4);
FULLADD_130: FULLADD port map (Sn1L3_14_Sn2L3_4,Sn1L3_14_Sn2L3_5,Sn1L3_14_Sn2L3_6,Sn1L4_14_Sn2L4_3,Sn1L4_15_Sn2L4_4);
FULLADD_131: FULLADD port map (Sn1L3_15_Sn2L3_4,Sn1L3_15_Sn2L3_5,Sn1L3_15_Sn2L3_6,Sn1L4_15_Sn2L4_3,Sn1L4_16_Sn2L4_4);
FULLADD_132: FULLADD port map (Sn1L3_16_Sn2L3_4,Sn1L3_16_Sn2L3_5,Sn1L3_16_Sn2L3_6,Sn1L4_16_Sn2L4_3,Sn1L4_17_Sn2L4_4);
FULLADD_133: FULLADD port map (Sn1L3_17_Sn2L3_4,Sn1L3_17_Sn2L3_5,Sn1L3_17_Sn2L3_6,Sn1L4_17_Sn2L4_3,Sn1L4_18_Sn2L4_4);
FULLADD_134: FULLADD port map (Sn1L3_18_Sn2L3_4,Sn1L3_18_Sn2L3_5,Sn1L3_18_Sn2L3_6,Sn1L4_18_Sn2L4_3,Sn1L4_19_Sn2L4_4);
FULLADD_135: FULLADD port map (Sn1L3_19_Sn2L3_4,Sn1L3_19_Sn2L3_5,Sn1L3_19_Sn2L3_6,Sn1L4_19_Sn2L4_3,Sn1L4_20_Sn2L4_4);
FULLADD_136: FULLADD port map (Sn1L3_20_Sn2L3_4,Sn1L3_20_Sn2L3_5,Sn1L3_20_Sn2L3_6,Sn1L4_20_Sn2L4_3,Sn1L4_21_Sn2L4_4);
FULLADD_137: FULLADD port map (Sn1L3_21_Sn2L3_4,Sn1L3_21_Sn2L3_5,Sn1L3_21_Sn2L3_6,Sn1L4_21_Sn2L4_3,Sn1L4_22_Sn2L4_4);
FULLADD_138: FULLADD port map (Sn1L3_22_Sn2L3_4,Sn1L3_22_Sn2L3_5,Sn1L3_22_Sn2L3_6,Sn1L4_22_Sn2L4_3,Sn1L4_23_Sn2L4_4);
FULLADD_139: FULLADD port map (Sn1L3_23_Sn2L3_4,Sn1L3_23_Sn2L3_5,Sn1L3_23_Sn2L3_6,Sn1L4_23_Sn2L4_3,Sn1L4_24_Sn2L4_4);
FULLADD_140: FULLADD port map (Sn1L3_24_Sn2L3_4,Sn1L3_24_Sn2L3_5,Sn1L3_24_Sn2L3_6,Sn1L4_24_Sn2L4_3,Sn1L4_25_Sn2L4_4);
FULLADD_141: FULLADD port map (Sn1L3_25_Sn2L3_4,A9B15,Sn1L3_25_Sn2L3_6,Sn1L4_25_Sn2L4_3,Sn1L4_26_Sn2L4_4);
FULLADD_142: FULLADD port map (Sn1L3_26_Sn2L3_4,A11B14,A10B15,Sn1L4_26_Sn2L4_3,Sn1L4_27_Sn2L4_4);
FULLADD_143: FULLADD port map (A13B13,A12B14,A11B15,Sn1L4_27_Sn2L4_3,Sn1L4_28_Sn2L4_4);

HALFADD_14: HALFADD port map (A3B0,A2B1,Sn1L5_4_Sn2L5_1,Sn1L5_5_Sn2L5_2);

FULLADD_144: FULLADD port map (Sn1L4_5_Sn2L4_1,A2B2,A1B3,Sn1L5_5_Sn2L5_1,Sn1L5_6_Sn2L5_2);
FULLADD_145: FULLADD port map (Sn1L4_6_Sn2L4_1,Sn1L4_6_Sn2L4_2,Sn1L4_6_Sn2L4_3,Sn1L5_6_Sn2L5_1,Sn1L5_7_Sn2L5_2);
FULLADD_146: FULLADD port map (Sn1L4_7_Sn2L4_1,Sn1L4_7_Sn2L4_2,Sn1L4_7_Sn2L4_3,Sn1L5_7_Sn2L5_1,Sn1L5_8_Sn2L5_2);
FULLADD_147: FULLADD port map (Sn1L4_8_Sn2L4_1,Sn1L4_8_Sn2L4_2,Sn1L4_8_Sn2L4_3,Sn1L5_8_Sn2L5_1,Sn1L5_9_Sn2L5_2);
FULLADD_148: FULLADD port map (Sn1L4_9_Sn2L4_1,Sn1L4_9_Sn2L4_2,Sn1L4_9_Sn2L4_3,Sn1L5_9_Sn2L5_1,Sn1L5_10_Sn2L5_2);
FULLADD_149: FULLADD port map (Sn1L4_10_Sn2L4_1,Sn1L4_10_Sn2L4_2,Sn1L4_10_Sn2L4_3,Sn1L5_10_Sn2L5_1,Sn1L5_11_Sn2L5_2);
FULLADD_150: FULLADD port map (Sn1L4_11_Sn2L4_1,Sn1L4_11_Sn2L4_2,Sn1L4_11_Sn2L4_3,Sn1L5_11_Sn2L5_1,Sn1L5_12_Sn2L5_2);
FULLADD_151: FULLADD port map (Sn1L4_12_Sn2L4_1,Sn1L4_12_Sn2L4_2,Sn1L4_12_Sn2L4_3,Sn1L5_12_Sn2L5_1,Sn1L5_13_Sn2L5_2);
FULLADD_152: FULLADD port map (Sn1L4_13_Sn2L4_1,Sn1L4_13_Sn2L4_2,Sn1L4_13_Sn2L4_3,Sn1L5_13_Sn2L5_1,Sn1L5_14_Sn2L5_2);
FULLADD_153: FULLADD port map (Sn1L4_14_Sn2L4_1,Sn1L4_14_Sn2L4_2,Sn1L4_14_Sn2L4_3,Sn1L5_14_Sn2L5_1,Sn1L5_15_Sn2L5_2);
FULLADD_154: FULLADD port map (Sn1L4_15_Sn2L4_1,Sn1L4_15_Sn2L4_2,Sn1L4_15_Sn2L4_3,Sn1L5_15_Sn2L5_1,Sn1L5_16_Sn2L5_2);
FULLADD_155: FULLADD port map (Sn1L4_16_Sn2L4_1,Sn1L4_16_Sn2L4_2,Sn1L4_16_Sn2L4_3,Sn1L5_16_Sn2L5_1,Sn1L5_17_Sn2L5_2);
FULLADD_156: FULLADD port map (Sn1L4_17_Sn2L4_1,Sn1L4_17_Sn2L4_2,Sn1L4_17_Sn2L4_3,Sn1L5_17_Sn2L5_1,Sn1L5_18_Sn2L5_2);
FULLADD_157: FULLADD port map (Sn1L4_18_Sn2L4_1,Sn1L4_18_Sn2L4_2,Sn1L4_18_Sn2L4_3,Sn1L5_18_Sn2L5_1,Sn1L5_19_Sn2L5_2);
FULLADD_158: FULLADD port map (Sn1L4_19_Sn2L4_1,Sn1L4_19_Sn2L4_2,Sn1L4_19_Sn2L4_3,Sn1L5_19_Sn2L5_1,Sn1L5_20_Sn2L5_2);
FULLADD_159: FULLADD port map (Sn1L4_20_Sn2L4_1,Sn1L4_20_Sn2L4_2,Sn1L4_20_Sn2L4_3,Sn1L5_20_Sn2L5_1,Sn1L5_21_Sn2L5_2);
FULLADD_160: FULLADD port map (Sn1L4_21_Sn2L4_1,Sn1L4_21_Sn2L4_2,Sn1L4_21_Sn2L4_3,Sn1L5_21_Sn2L5_1,Sn1L5_22_Sn2L5_2);
FULLADD_161: FULLADD port map (Sn1L4_22_Sn2L4_1,Sn1L4_22_Sn2L4_2,Sn1L4_22_Sn2L4_3,Sn1L5_22_Sn2L5_1,Sn1L5_23_Sn2L5_2);
FULLADD_162: FULLADD port map (Sn1L4_23_Sn2L4_1,Sn1L4_23_Sn2L4_2,Sn1L4_23_Sn2L4_3,Sn1L5_23_Sn2L5_1,Sn1L5_24_Sn2L5_2);
FULLADD_163: FULLADD port map (Sn1L4_24_Sn2L4_1,Sn1L4_24_Sn2L4_2,Sn1L4_24_Sn2L4_3,Sn1L5_24_Sn2L5_1,Sn1L5_25_Sn2L5_2);
FULLADD_164: FULLADD port map (Sn1L4_25_Sn2L4_1,Sn1L4_25_Sn2L4_2,Sn1L4_25_Sn2L4_3,Sn1L5_25_Sn2L5_1,Sn1L5_26_Sn2L5_2);
FULLADD_165: FULLADD port map (Sn1L4_26_Sn2L4_1,Sn1L4_26_Sn2L4_2,Sn1L4_26_Sn2L4_3,Sn1L5_26_Sn2L5_1,Sn1L5_27_Sn2L5_2);
FULLADD_166: FULLADD port map (Sn1L4_27_Sn2L4_1,Sn1L4_27_Sn2L4_2,Sn1L4_27_Sn2L4_3,Sn1L5_27_Sn2L5_1,Sn1L5_28_Sn2L5_2);
FULLADD_167: FULLADD port map (Sn1L4_28_Sn2L4_1,Sn1L4_28_Sn2L4_2,A12B15,Sn1L5_28_Sn2L5_1,Sn1L5_29_Sn2L5_2);
FULLADD_168: FULLADD port map (A15B13,Sn1L4_29_Sn2L4_2,A14B14,Sn1L5_29_Sn2L5_1,Sn1L5_30_Sn2L5_2);

HALFADD_15: HALFADD port map (A2B0,A1B1,Sn1L6_3_Sn2L6_1,Sn1L6_4_Sn2L6_2);

FULLADD_169: FULLADD port map (Sn1L5_4_Sn2L5_1,A1B2,A0B3,Sn1L6_4_Sn2L6_1,Sn1L6_5_Sn2L6_2);
FULLADD_170: FULLADD port map (Sn1L5_5_Sn2L5_1,Sn1L5_5_Sn2L5_2,A0B4,Sn1L6_5_Sn2L6_1,Sn1L6_6_Sn2L6_2);
FULLADD_171: FULLADD port map (Sn1L5_6_Sn2L5_1,Sn1L5_6_Sn2L5_2,A0B5,Sn1L6_6_Sn2L6_1,Sn1L6_7_Sn2L6_2);
FULLADD_172: FULLADD port map (Sn1L5_7_Sn2L5_1,Sn1L5_7_Sn2L5_2,Sn1L4_7_Sn2L4_4,Sn1L6_7_Sn2L6_1,Sn1L6_8_Sn2L6_2);
FULLADD_173: FULLADD port map (Sn1L5_8_Sn2L5_1,Sn1L5_8_Sn2L5_2,Sn1L4_8_Sn2L4_4,Sn1L6_8_Sn2L6_1,Sn1L6_9_Sn2L6_2);
FULLADD_174: FULLADD port map (Sn1L5_9_Sn2L5_1,Sn1L5_9_Sn2L5_2,Sn1L4_9_Sn2L4_4,Sn1L6_9_Sn2L6_1,Sn1L6_10_Sn2L6_2);
FULLADD_175: FULLADD port map (Sn1L5_10_Sn2L5_1,Sn1L5_10_Sn2L5_2,Sn1L4_10_Sn2L4_4,Sn1L6_10_Sn2L6_1,Sn1L6_11_Sn2L6_2);
FULLADD_176: FULLADD port map (Sn1L5_11_Sn2L5_1,Sn1L5_11_Sn2L5_2,Sn1L4_11_Sn2L4_4,Sn1L6_11_Sn2L6_1,Sn1L6_12_Sn2L6_2);
FULLADD_177: FULLADD port map (Sn1L5_12_Sn2L5_1,Sn1L5_12_Sn2L5_2,Sn1L4_12_Sn2L4_4,Sn1L6_12_Sn2L6_1,Sn1L6_13_Sn2L6_2);
FULLADD_178: FULLADD port map (Sn1L5_13_Sn2L5_1,Sn1L5_13_Sn2L5_2,Sn1L4_13_Sn2L4_4,Sn1L6_13_Sn2L6_1,Sn1L6_14_Sn2L6_2);
FULLADD_179: FULLADD port map (Sn1L5_14_Sn2L5_1,Sn1L5_14_Sn2L5_2,Sn1L4_14_Sn2L4_4,Sn1L6_14_Sn2L6_1,Sn1L6_15_Sn2L6_2);
FULLADD_180: FULLADD port map (Sn1L5_15_Sn2L5_1,Sn1L5_15_Sn2L5_2,Sn1L4_15_Sn2L4_4,Sn1L6_15_Sn2L6_1,Sn1L6_16_Sn2L6_2);
FULLADD_181: FULLADD port map (Sn1L5_16_Sn2L5_1,Sn1L5_16_Sn2L5_2,Sn1L4_16_Sn2L4_4,Sn1L6_16_Sn2L6_1,Sn1L6_17_Sn2L6_2);
FULLADD_182: FULLADD port map (Sn1L5_17_Sn2L5_1,Sn1L5_17_Sn2L5_2,Sn1L4_17_Sn2L4_4,Sn1L6_17_Sn2L6_1,Sn1L6_18_Sn2L6_2);
FULLADD_183: FULLADD port map (Sn1L5_18_Sn2L5_1,Sn1L5_18_Sn2L5_2,Sn1L4_18_Sn2L4_4,Sn1L6_18_Sn2L6_1,Sn1L6_19_Sn2L6_2);
FULLADD_184: FULLADD port map (Sn1L5_19_Sn2L5_1,Sn1L5_19_Sn2L5_2,Sn1L4_19_Sn2L4_4,Sn1L6_19_Sn2L6_1,Sn1L6_20_Sn2L6_2);
FULLADD_185: FULLADD port map (Sn1L5_20_Sn2L5_1,Sn1L5_20_Sn2L5_2,Sn1L4_20_Sn2L4_4,Sn1L6_20_Sn2L6_1,Sn1L6_21_Sn2L6_2);
FULLADD_186: FULLADD port map (Sn1L5_21_Sn2L5_1,Sn1L5_21_Sn2L5_2,Sn1L4_21_Sn2L4_4,Sn1L6_21_Sn2L6_1,Sn1L6_22_Sn2L6_2);
FULLADD_187: FULLADD port map (Sn1L5_22_Sn2L5_1,Sn1L5_22_Sn2L5_2,Sn1L4_22_Sn2L4_4,Sn1L6_22_Sn2L6_1,Sn1L6_23_Sn2L6_2);
FULLADD_188: FULLADD port map (Sn1L5_23_Sn2L5_1,Sn1L5_23_Sn2L5_2,Sn1L4_23_Sn2L4_4,Sn1L6_23_Sn2L6_1,Sn1L6_24_Sn2L6_2);
FULLADD_189: FULLADD port map (Sn1L5_24_Sn2L5_1,Sn1L5_24_Sn2L5_2,Sn1L4_24_Sn2L4_4,Sn1L6_24_Sn2L6_1,Sn1L6_25_Sn2L6_2);
FULLADD_190: FULLADD port map (Sn1L5_25_Sn2L5_1,Sn1L5_25_Sn2L5_2,Sn1L4_25_Sn2L4_4,Sn1L6_25_Sn2L6_1,Sn1L6_26_Sn2L6_2);
FULLADD_191: FULLADD port map (Sn1L5_26_Sn2L5_1,Sn1L5_26_Sn2L5_2,Sn1L4_26_Sn2L4_4,Sn1L6_26_Sn2L6_1,Sn1L6_27_Sn2L6_2);
FULLADD_192: FULLADD port map (Sn1L5_27_Sn2L5_1,Sn1L5_27_Sn2L5_2,Sn1L4_27_Sn2L4_4,Sn1L6_27_Sn2L6_1,Sn1L6_28_Sn2L6_2);
FULLADD_193: FULLADD port map (Sn1L5_28_Sn2L5_1,Sn1L5_28_Sn2L5_2,Sn1L4_28_Sn2L4_4,Sn1L6_28_Sn2L6_1,Sn1L6_29_Sn2L6_2);
FULLADD_194: FULLADD port map (Sn1L5_29_Sn2L5_1,Sn1L5_29_Sn2L5_2,A13B15,Sn1L6_29_Sn2L6_1,Sn1L6_30_Sn2L6_2);
FULLADD_195: FULLADD port map (A15B14,Sn1L5_30_Sn2L5_2,A14B15,Sn1L6_30_Sn2L6_1,Sn1L6_31_Sn2L6_2);

Ain <= '0' & A15B15 & Sn1L6_30_Sn2L6_1 & Sn1L6_29_Sn2L6_1 & Sn1L6_28_Sn2L6_1 & Sn1L6_27_Sn2L6_1 & Sn1L6_26_Sn2L6_1 & Sn1L6_25_Sn2L6_1 & Sn1L6_24_Sn2L6_1 & Sn1L6_23_Sn2L6_1 & Sn1L6_22_Sn2L6_1 & Sn1L6_21_Sn2L6_1 & Sn1L6_20_Sn2L6_1 & Sn1L6_19_Sn2L6_1 & Sn1L6_18_Sn2L6_1 & Sn1L6_17_Sn2L6_1 & Sn1L6_16_Sn2L6_1 & Sn1L6_15_Sn2L6_1 & Sn1L6_14_Sn2L6_1 & Sn1L6_13_Sn2L6_1 & Sn1L6_12_Sn2L6_1 & Sn1L6_11_Sn2L6_1 & Sn1L6_10_Sn2L6_1 & Sn1L6_9_Sn2L6_1 & Sn1L6_8_Sn2L6_1 & Sn1L6_7_Sn2L6_1 & Sn1L6_6_Sn2L6_1 & Sn1L6_5_Sn2L6_1 & Sn1L6_4_Sn2L6_1 &  Sn1L6_3_Sn2L6_1 & A1B0 & A0B0;
Bin <= '0' & Sn1L6_31_Sn2L6_2 & Sn1L6_30_Sn2L6_2 & Sn1L6_29_Sn2L6_2 & Sn1L6_28_Sn2L6_2 & Sn1L6_27_Sn2L6_2 & Sn1L6_26_Sn2L6_2 & Sn1L6_25_Sn2L6_2 & Sn1L6_24_Sn2L6_2 & Sn1L6_23_Sn2L6_2 & Sn1L6_22_Sn2L6_2 & Sn1L6_21_Sn2L6_2 & Sn1L6_20_Sn2L6_2 & Sn1L6_19_Sn2L6_2 & Sn1L6_18_Sn2L6_2 & Sn1L6_17_Sn2L6_2 & Sn1L6_16_Sn2L6_2 & Sn1L6_15_Sn2L6_2 & Sn1L6_14_Sn2L6_2 & Sn1L6_13_Sn2L6_2 & Sn1L6_12_Sn2L6_2 & Sn1L6_11_Sn2L6_2 & Sn1L6_10_Sn2L6_2 & Sn1L6_9_Sn2L6_2 & Sn1L6_8_Sn2L6_2 & Sn1L6_7_Sn2L6_2 & Sn1L6_6_Sn2L6_2 & Sn1L6_5_Sn2L6_2 & Sn1L6_4_Sn2L6_2 &  A0B2 & A0B1 & '0';

ADD: brentkung_32bit_adder port map(Ain,Bin,'0',M,nocarry);

END a1;